*TB_SUN_TR_SKY130NM/TB_NCM

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc 0 pwl 0 0 10n {AVDD}



VIN VIN 0 dc 0 sin (0 10m 1G 1u 0 0 )

*- Make a bias source
R1 VDD_1V8 VBIAS 10k
XM1 VBIAS VBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=0.2 W=1
R2 VBIAS VG 100k

*- Common source amplifier
C1 VIN VG 1p
R3 VDD_1V8 VOUT 5k
XM2 VOUT VG VSS VSS sky130_fd_pr__nfet_01v8 L=0.2 W=1 M=10

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0
tran 10p 1.1u 1.09u
write
quit

.endc

.end
